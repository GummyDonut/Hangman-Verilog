library verilog;
use verilog.vl_types.all;
entity storageFinal_vlg_sample_tst is
    port(
        \Clock\         : in     vl_logic;
        Resetn          : in     vl_logic;
        clock           : in     vl_logic;
        confirm         : in     vl_logic;
        up_down         : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end storageFinal_vlg_sample_tst;
