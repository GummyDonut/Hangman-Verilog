library verilog;
use verilog.vl_types.all;
entity statemachineforpigs_vlg_check_tst is
    port(
        T               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end statemachineforpigs_vlg_check_tst;
