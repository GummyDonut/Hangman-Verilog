library verilog;
use verilog.vl_types.all;
entity statemachineforpigs_vlg_vec_tst is
end statemachineforpigs_vlg_vec_tst;
