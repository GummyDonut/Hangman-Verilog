library verilog;
use verilog.vl_types.all;
entity storageFinal_vlg_vec_tst is
end storageFinal_vlg_vec_tst;
